module XilinxU250Board (
    input pcie_mgt_clkn,
    input pcie_mgt_clkp,
    input pcie_perstn_rst,
    input  [15:0] pci_exp_rxn,
    input  [15:0] pci_exp_rxp,
    output [15:0] pci_exp_txn,
    output [15:0] pci_exp_txp
);

wire sys_clk;
wire sys_clk_gt;
wire axi_aclk;
wire axi_aresetn;

wire [63:0] m_axi_awaddr;
wire [7:0] m_axi_awlen;
wire [2:0] m_axi_awsize;
wire [1:0] m_axi_awburst;
wire m_axi_awlock;
wire [3:0] m_axi_awcache;
wire [2:0] m_axi_awprot;
wire m_axi_awvalid;
wire m_axi_awready;
wire [511:0] m_axi_wdata;
wire [63:0] m_axi_wstrb;
wire m_axi_wlast;
wire m_axi_wvalid;
wire m_axi_wready;
wire [1:0] m_axi_bresp;
wire m_axi_bvalid;
wire m_axi_bready;
wire [63:0] m_axi_araddr;
wire [7:0] m_axi_arlen;
wire [2:0] m_axi_arsize;
wire [1:0] m_axi_arburst;
wire m_axi_arlock;
wire [3:0] m_axi_arcache;
wire [2:0] m_axi_arprot;
wire m_axi_arvalid;
wire m_axi_arready;
wire [511:0] m_axi_rdata;
wire [1:0] m_axi_rresp;
wire m_axi_rlast;
wire m_axi_rvalid;
wire m_axi_rready;

wire bram_rst_a;
wire bram_clk_a;
wire bram_en_a;
wire [63:0] bram_we_a;
wire [18:0] bram_addr_a;
wire [511:0] bram_wrdata_a;
wire [511:0] bram_rddata_a;
wire bram_rst_b;
wire bram_clk_b;
wire bram_en_b;
wire [63:0] bram_we_b;
wire [18:0] bram_addr_b;
wire [511:0] bram_wrdata_b;
wire [511:0] bram_rddata_b;

wire [31:0] m_axil_awaddr;
wire [2:0] m_axil_awprot;
wire m_axil_awvalid;
wire m_axil_awready;
wire [31:0] m_axil_wdata;
wire [3:0] m_axil_wstrb;
wire m_axil_wvalid;
wire m_axil_wready;
wire m_axil_bvalid;
wire [1:0] m_axil_bresp;
wire m_axil_bready;
wire [31:0] m_axil_araddr;
wire [2:0] m_axil_arprot;
wire m_axil_arvalid;
wire m_axil_arready;
wire [31:0] m_axil_rdata;
wire [1:0] m_axil_rresp;
wire m_axil_rvalid;
wire m_axil_rready;

wire bram_rst_a_0;
wire bram_clk_a_0;
wire bram_en_a_0;
wire [3:0] bram_we_a_0;
wire [14:0] bram_addr_a_0;
wire [31:0] bram_wrdata_a_0;
wire [31:0] bram_rddata_a_0;
wire bram_rst_b_0;
wire bram_clk_b_0;
wire bram_en_b_0;
wire [3:0] bram_we_b_0;
wire [14:0] bram_addr_b_0;
wire [31:0] bram_wrdata_b_0;
wire [31:0] bram_rddata_b_0;

IBUFDS_GTE4 #(
  .REFCLK_HROW_CK_SEL(2'b00)
)
IBUFDS_inst (
   .O(sys_clk_gt),         // 1-bit output: Refer to Transceiver User Guide.
   .I (pcie_mgt_clkp),     // 1-bit input: Refer to Transceiver User Guide.
   .IB(pcie_mgt_clkn),      // 1-bit input: Refer to Transceiver User Guide.
   .CEB(1'b0),
   .ODIV2(sys_clk)
);

xdma_0 xdma_0 (
  .sys_clk(sys_clk),                                    // input wire sys_clk
  .sys_clk_gt(sys_clk_gt),                                 // input wire sys_clk_gt
  .sys_rst_n(pcie_perstn_rst),                          // input wire sys_rst_n
  .user_lnk_up(),                                       // output wire user_lnk_up
  .pci_exp_txp(pci_exp_txp),                            // output wire [15 : 0] pci_exp_txp
  .pci_exp_txn(pci_exp_txn),                            // output wire [15 : 0] pci_exp_txn
  .pci_exp_rxp(pci_exp_rxp),                            // input wire [15 : 0] pci_exp_rxp
  .pci_exp_rxn(pci_exp_rxn),                            // input wire [15 : 0] pci_exp_rxn
  .axi_aclk(axi_aclk),                                  // output wire axi_aclk
  .axi_aresetn(axi_aresetn),                            // output wire axi_aresetn
  .usr_irq_req(1'b0),                                   // input wire [0 : 0] usr_irq_req
  .usr_irq_ack(),                                       // output wire [0 : 0] usr_irq_ack
  .msi_enable(),                                        // output wire msi_enable
  .msi_vector_width(),                                  // output wire [2 : 0] msi_vector_width

  .m_axi_awready(m_axi_awready),                        // input wire m_axi_awready
  .m_axi_wready(m_axi_wready),                          // input wire m_axi_wready
  .m_axi_bid(4'b0),                                // input wire [3 : 0] m_axi_bid
  .m_axi_bresp(m_axi_bresp),                            // input wire [1 : 0] m_axi_bresp
  .m_axi_bvalid(m_axi_bvalid),                          // input wire m_axi_bvalid
  .m_axi_arready(m_axi_arready),                        // input wire m_axi_arready
  .m_axi_rid(4'b0),                                // input wire [3 : 0] m_axi_rid
  .m_axi_rdata(m_axi_rdata),                            // input wire [511 : 0] m_axi_rdata
  .m_axi_rresp(m_axi_rresp),                            // input wire [1 : 0] m_axi_rresp
  .m_axi_rlast(m_axi_rlast),                            // input wire m_axi_rlast
  .m_axi_rvalid(m_axi_rvalid),                          // input wire m_axi_rvalid
  .m_axi_awid(),                              // output wire [3 : 0] m_axi_awid
  .m_axi_awaddr(m_axi_awaddr),                          // output wire [63 : 0] m_axi_awaddr
  .m_axi_awlen(m_axi_awlen),                            // output wire [7 : 0] m_axi_awlen
  .m_axi_awsize(m_axi_awsize),                          // output wire [2 : 0] m_axi_awsize
  .m_axi_awburst(m_axi_awburst),                        // output wire [1 : 0] m_axi_awburst
  .m_axi_awprot(m_axi_awprot),                          // output wire [2 : 0] m_axi_awprot
  .m_axi_awvalid(m_axi_awvalid),                        // output wire m_axi_awvalid
  .m_axi_awlock(m_axi_awlock),                          // output wire m_axi_awlock
  .m_axi_awcache(m_axi_awcache),                        // output wire [3 : 0] m_axi_awcache
  .m_axi_wdata(m_axi_wdata),                            // output wire [511 : 0] m_axi_wdata
  .m_axi_wstrb(m_axi_wstrb),                            // output wire [63 : 0] m_axi_wstrb
  .m_axi_wlast(m_axi_wlast),                            // output wire m_axi_wlast
  .m_axi_wvalid(m_axi_wvalid),                          // output wire m_axi_wvalid
  .m_axi_bready(m_axi_bready),                          // output wire m_axi_bready
  .m_axi_arid(),                              // output wire [3 : 0] m_axi_arid
  .m_axi_araddr(m_axi_araddr),                          // output wire [63 : 0] m_axi_araddr
  .m_axi_arlen(m_axi_arlen),                            // output wire [7 : 0] m_axi_arlen
  .m_axi_arsize(m_axi_arsize),                          // output wire [2 : 0] m_axi_arsize
  .m_axi_arburst(m_axi_arburst),                        // output wire [1 : 0] m_axi_arburst
  .m_axi_arprot(m_axi_arprot),                          // output wire [2 : 0] m_axi_arprot
  .m_axi_arvalid(m_axi_arvalid),                        // output wire m_axi_arvalid
  .m_axi_arlock(m_axi_arlock),                          // output wire m_axi_arlock
  .m_axi_arcache(m_axi_arcache),                        // output wire [3 : 0] m_axi_arcache
  .m_axi_rready(m_axi_rready),                          // output wire m_axi_rready

  .m_axil_awaddr(m_axil_awaddr),                        // output wire [31 : 0] m_axil_awaddr
  .m_axil_awprot(m_axil_awprot),                        // output wire [2 : 0] m_axil_awprot
  .m_axil_awvalid(m_axil_awvalid),                      // output wire m_axil_awvalid
  .m_axil_awready(m_axil_awready),                      // input wire m_axil_awready
  .m_axil_wdata(m_axil_wdata),                          // output wire [31 : 0] m_axil_wdata
  .m_axil_wstrb(m_axil_wstrb),                          // output wire [3 : 0] m_axil_wstrb
  .m_axil_wvalid(m_axil_wvalid),                        // output wire m_axil_wvalid
  .m_axil_wready(m_axil_wready),                        // input wire m_axil_wready
  .m_axil_bvalid(m_axil_bvalid),                        // input wire m_axil_bvalid
  .m_axil_bresp(m_axil_bresp),                          // input wire [1 : 0] m_axil_bresp
  .m_axil_bready(m_axil_bready),                        // output wire m_axil_bready
  .m_axil_araddr(m_axil_araddr),                        // output wire [31 : 0] m_axil_araddr
  .m_axil_arprot(m_axil_arprot),                        // output wire [2 : 0] m_axil_arprot
  .m_axil_arvalid(m_axil_arvalid),                      // output wire m_axil_arvalid
  .m_axil_arready(m_axil_arready),                      // input wire m_axil_arready
  .m_axil_rdata(m_axil_rdata),                          // input wire [31 : 0] m_axil_rdata
  .m_axil_rresp(m_axil_rresp),                          // input wire [1 : 0] m_axil_rresp
  .m_axil_rvalid(m_axil_rvalid),                        // input wire m_axil_rvalid
  .m_axil_rready(m_axil_rready),                        // output wire m_axil_rready
  .cfg_mgmt_addr(),                                     // input wire [18 : 0] cfg_mgmt_addr
  .cfg_mgmt_write(),                                    // input wire cfg_mgmt_write
  .cfg_mgmt_write_data(),                               // input wire [31 : 0] cfg_mgmt_write_data
  .cfg_mgmt_byte_enable(),                              // input wire [3 : 0] cfg_mgmt_byte_enable
  .cfg_mgmt_read(),                                     // input wire cfg_mgmt_read
  .cfg_mgmt_read_data(),                                // output wire [31 : 0] cfg_mgmt_read_data
  .cfg_mgmt_read_write_done()                           // output wire cfg_mgmt_read_write_done
);

ila_0 xdma_dma_ila (
  .clk(axi_aclk), // input wire clk
  .probe0 (m_axi_wready), // input wire [0:0] probe0  
  .probe1 (m_axi_awaddr), // input wire [63:0]  probe1 
  .probe2 (m_axi_bresp), // input wire [1:0]  probe2 
  .probe3 (m_axi_bvalid), // input wire [0:0]  probe3 
  .probe4 (m_axi_bready), // input wire [0:0]  probe4 
  .probe5 (m_axi_araddr), // input wire [63:0]  probe5 
  .probe6 (m_axi_rready), // input wire [0:0]  probe6 
  .probe7 (m_axi_wvalid), // input wire [0:0]  probe7 
  .probe8 (m_axi_arvalid), // input wire [0:0]  probe8 
  .probe9 (m_axi_arready), // input wire [0:0]  probe9 
  .probe10(m_axi_rdata), // input wire [511:0]  probe10 
  .probe11(m_axi_awvalid), // input wire [0:0]  probe11 
  .probe12(m_axi_awready), // input wire [0:0]  probe12 
  .probe13(m_axi_rresp), // input wire [1:0]  probe13 
  .probe14(m_axi_wdata), // input wire [511:0]  probe14 
  .probe15(m_axi_wstrb), // input wire [63:0]  probe15 
  .probe16(m_axi_rvalid), // input wire [0:0]  probe16 
  .probe17(m_axi_arprot), // input wire [2:0]  probe17 
  .probe18(m_axi_awprot), // input wire [2:0]  probe18 
  .probe19(1'b0), // input wire [0:0]  probe19 
  .probe20(1'b0), // input wire [0:0]  probe20 
  .probe21(m_axi_awlen), // input wire [7:0]  probe21 
  .probe22(1'b0), // input wire [0:0]  probe22 
  .probe23(m_axi_awsize), // input wire [2:0]  probe23 
  .probe24(m_axi_awburst), // input wire [1:0]  probe24 
  .probe25(4'b0), // input wire [0:0]  probe25 
  .probe26(m_axi_awlock), // input wire [0:0]  probe26 
  .probe27(m_axi_arlen), // input wire [7:0]  probe27 
  .probe28(m_axi_arsize), // input wire [2:0]  probe28 
  .probe29(m_axi_arburst), // input wire [1:0]  probe29 
  .probe30(m_axi_arlock), // input wire [0:0]  probe30 
  .probe31(m_axi_arcache), // input wire [3:0]  probe31 
  .probe32(m_axi_awcache), // input wire [3:0]  probe32 
  .probe33(4'b0), // input wire [3:0]  probe33 
  .probe34(3'b0), // input wire [3:0]  probe34 
  .probe35(1'b0), // input wire [0:0]  probe35 
  .probe36(4'b0), // input wire [3:0]  probe36 
  .probe37(4'b0), // input wire [3:0]  probe37 
  .probe38(1'b0), // input wire [0:0]  probe38 
  .probe39(1'b0), // input wire [0:0]  probe39 
  .probe40(1'b0), // input wire [0:0]  probe40 
  .probe41(m_axi_rlast), // input wire [0:0]  probe41 
  .probe42(1'b0), // input wire [0:0]  probe42  
  .probe43(m_axi_wlast) // input wire [0:0]  probe43
);

axi_bram_ctrl_0_512 axi_bram_ctrl_0_512 (
  .s_axi_aclk(axi_aclk),        // input wire s_axi_aclk
  .s_axi_aresetn(axi_aresetn),  // input wire s_axi_aresetn
  .s_axi_awaddr(m_axi_awaddr),    // input wire [18 : 0] s_axi_awaddr
  .s_axi_awlen(m_axi_awlen),      // input wire [7 : 0] s_axi_awlen
  .s_axi_awsize(m_axi_awsize),    // input wire [2 : 0] s_axi_awsize
  .s_axi_awburst(m_axi_awburst),  // input wire [1 : 0] s_axi_awburst
  .s_axi_awlock(m_axi_awlock),    // input wire s_axi_awlock
  .s_axi_awcache(m_axi_awcache),  // input wire [3 : 0] s_axi_awcache
  .s_axi_awprot(m_axi_awprot),    // input wire [2 : 0] s_axi_awprot
  .s_axi_awvalid(m_axi_awvalid),  // input wire s_axi_awvalid
  .s_axi_awready(m_axi_awready),  // output wire s_axi_awready
  .s_axi_wdata(m_axi_wdata),      // input wire [511 : 0] s_axi_wdata
  .s_axi_wstrb(m_axi_wstrb),      // input wire [63 : 0] s_axi_wstrb
  .s_axi_wlast(m_axi_wlast),      // input wire s_axi_wlast
  .s_axi_wvalid(m_axi_wvalid),    // input wire s_axi_wvalid
  .s_axi_wready(m_axi_wready),    // output wire s_axi_wready
  .s_axi_bresp(m_axi_bresp),      // output wire [1 : 0] s_axi_bresp
  .s_axi_bvalid(m_axi_bvalid),    // output wire s_axi_bvalid
  .s_axi_bready(m_axi_bready),    // input wire s_axi_bready
  .s_axi_araddr(m_axi_araddr),    // input wire [18 : 0] s_axi_araddr
  .s_axi_arlen(m_axi_arlen),      // input wire [7 : 0] s_axi_arlen
  .s_axi_arsize(m_axi_arsize),    // input wire [2 : 0] s_axi_arsize
  .s_axi_arburst(m_axi_arburst),  // input wire [1 : 0] s_axi_arburst
  .s_axi_arlock(m_axi_arlock),    // input wire s_axi_arlock
  .s_axi_arcache(m_axi_arcache),  // input wire [3 : 0] s_axi_arcache
  .s_axi_arprot(m_axi_arprot),    // input wire [2 : 0] s_axi_arprot
  .s_axi_arvalid(m_axi_arvalid),  // input wire s_axi_arvalid
  .s_axi_arready(m_axi_arready),  // output wire s_axi_arready
  .s_axi_rdata(m_axi_rdata),      // output wire [511 : 0] s_axi_rdata
  .s_axi_rresp(m_axi_rresp),      // output wire [1 : 0] s_axi_rresp
  .s_axi_rlast(m_axi_rlast),      // output wire s_axi_rlast
  .s_axi_rvalid(m_axi_rvalid),    // output wire s_axi_rvalid
  .s_axi_rready(m_axi_rready),    // input wire s_axi_rready
  .bram_rst_a(bram_rst_a),        // output wire bram_rst_a
  .bram_clk_a(bram_clk_a),        // output wire bram_clk_a
  .bram_en_a(bram_en_a),          // output wire bram_en_a
  .bram_we_a(bram_we_a),          // output wire [63 : 0] bram_we_a
  .bram_addr_a(bram_addr_a),      // output wire [18 : 0] bram_addr_a
  .bram_wrdata_a(bram_wrdata_a),  // output wire [511 : 0] bram_wrdata_a
  .bram_rddata_a(bram_rddata_a),  // input wire [511 : 0] bram_rddata_a
  .bram_rst_b(bram_rst_b),        // output wire bram_rst_b
  .bram_clk_b(bram_clk_b),        // output wire bram_clk_b
  .bram_en_b(bram_en_b),          // output wire bram_en_b
  .bram_we_b(bram_we_b),          // output wire [63 : 0] bram_we_b
  .bram_addr_b(bram_addr_b),      // output wire [18 : 0] bram_addr_b
  .bram_wrdata_b(bram_wrdata_b),  // output wire [511 : 0] bram_wrdata_b
  .bram_rddata_b(bram_rddata_b)  // input wire [511 : 0] bram_rddata_b
);

bram_0_512 bram_0_512 (
  .clka(bram_clk_a),       // input wire clka
  .ena(bram_en_a),         // input wire ena
  .wea(bram_we_a),         // input wire [0 : 0] wea
  .addra(bram_addr_a),     // input wire [9 : 0] addra
  .dina(bram_wrdata_a),    // input wire [511 : 0] dina
  .douta(bram_rddata_a),   // output wire [511 : 0] douta
  .clkb(bram_clk_b),       // input wire clkb
  .enb(bram_en_b),         // input wire enb
  .web(bram_we_b),         // input wire [0 : 0] web
  .addrb(bram_addr_b),     // input wire [9 : 0] addrb
  .dinb(bram_wrdata_b),    // input wire [511 : 0] dinb
  .doutb(bram_rddata_b)    // output wire [511 : 0] doutb
);

axi_lite_bram_ctrl_0_32 axi_lite_bram_ctrl_0_32 (
  .s_axi_aclk(axi_aclk),            // input wire s_axi_aclk
  .s_axi_aresetn(axi_aresetn),      // input wire s_axi_aresetn
  .s_axi_awaddr(m_axil_awaddr),     // input wire [14 : 0] s_axi_awaddr
  .s_axi_awprot(m_axil_awprot),     // input wire [2 : 0] s_axi_awprot
  .s_axi_awvalid(m_axil_awvalid),   // input wire s_axi_awvalid
  .s_axi_awready(m_axil_awready),   // output wire s_axi_awready
  .s_axi_wdata(m_axil_wdata),       // input wire [31 : 0] s_axi_wdata
  .s_axi_wstrb(m_axil_wstrb),       // input wire [3 : 0] s_axi_wstrb
  .s_axi_wvalid(m_axil_wvalid),     // input wire s_axi_wvalid
  .s_axi_wready(m_axil_wready),     // output wire s_axi_wready
  .s_axi_bresp(m_axil_bresp),       // output wire [1 : 0] s_axi_bresp
  .s_axi_bvalid(m_axil_bvalid),     // output wire s_axi_bvalid
  .s_axi_bready(m_axil_bready),     // input wire s_axi_bready
  .s_axi_araddr(m_axil_araddr),     // input wire [14 : 0] s_axi_araddr
  .s_axi_arprot(m_axil_arprot),     // input wire [2 : 0] s_axi_arprot
  .s_axi_arvalid(m_axil_arvalid),   // input wire s_axi_arvalid
  .s_axi_arready(m_axil_arready),   // output wire s_axi_arready
  .s_axi_rdata(m_axil_rdata),       // output wire [31 : 0] s_axi_rdata
  .s_axi_rresp(m_axil_rresp),       // output wire [1 : 0] s_axi_rresp
  .s_axi_rvalid(m_axil_rvalid),     // output wire s_axi_rvalid
  .s_axi_rready(m_axil_rready),     // input wire s_axi_rready
  .bram_rst_a(bram_rst_a_0),        // output wire bram_rst_a
  .bram_clk_a(bram_clk_a_0),        // output wire bram_clk_a
  .bram_en_a(bram_en_a_0),          // output wire bram_en_a
  .bram_we_a(bram_we_a_0),          // output wire [3 : 0] bram_we_a
  .bram_addr_a(bram_addr_a_0),      // output wire [14 : 0] bram_addr_a
  .bram_wrdata_a(bram_wrdata_a_0),  // output wire [31 : 0] bram_wrdata_a
  .bram_rddata_a(bram_rddata_a_0),  // input wire [31 : 0] bram_rddata_a
  .bram_rst_b(bram_rst_b_0),        // output wire bram_rst_b
  .bram_clk_b(bram_clk_b_0),        // output wire bram_clk_b
  .bram_en_b(bram_en_b_0),          // output wire bram_en_b
  .bram_we_b(bram_we_b_0),          // output wire [3 : 0] bram_we_b
  .bram_addr_b(bram_addr_b_0),      // output wire [14 : 0] bram_addr_b
  .bram_wrdata_b(bram_wrdata_b_0),  // output wire [31 : 0] bram_wrdata_b
  .bram_rddata_b(bram_rddata_b_0)   // input wire [31 : 0] bram_rddata_b
);

bram_0_32 bram_0_32 (
  .clka(bram_clk_a_0),       // input wire clka
  .ena(bram_en_a_0),         // input wire ena
  .wea(bram_we_a_0),         // input wire [0 : 0] wea
  .addra(bram_addr_a_0),     // input wire [9 : 0] addra
  .dina(bram_wrdata_a_0),    // input wire [31 : 0] dina
  .douta(bram_rddata_a_0),   // output wire [31 : 0] douta
  .clkb(bram_clk_b_0),       // input wire clkb
  .enb(bram_en_b_0),         // input wire enb
  .web(bram_we_b_0),         // input wire [0 : 0] web
  .addrb(bram_addr_b_0),     // input wire [9 : 0] addrb
  .dinb(bram_wrdata_b_0),    // input wire [31 : 0] dinb
  .doutb(bram_rddata_b_0)    // output wire [31 : 0] doutb
);

ila_0 xdma_mmio_ila (
  .clk    (axi_aclk), // input wire clk
  .probe0(axi_aresetn),      // input wire s_axi_aresetn
  .probe1(m_axil_awaddr),     // input wire [14 : 0] s_axi_awaddr
  .probe2(m_axil_awprot),     // input wire [2 : 0] s_axi_awprot
  .probe3(m_axil_awvalid),   // input wire s_axi_awvalid
  .probe4(m_axil_awready),   // output wire s_axi_awready
  .probe5(m_axil_wdata),       // input wire [31 : 0] s_axi_wdata
  .probe6(m_axil_wstrb),       // input wire [3 : 0] s_axi_wstrb
  .probe7(m_axil_wvalid),     // input wire s_axi_wvalid
  .probe8(m_axil_wready),     // output wire s_axi_wready
  .probe9(m_axil_bresp),       // output wire [1 : 0] s_axi_bresp
  .probe10(m_axil_bvalid),     // output wire s_axi_bvalid
  .probe11(m_axil_bready),     // input wire s_axi_bready
  .probe12(m_axil_araddr),     // input wire [14 : 0] s_axi_araddr
  .probe13(m_axil_arprot),     // input wire [2 : 0] s_axi_arprot
  .probe14(m_axil_arvalid),   // input wire s_axi_arvalid
  .probe15(m_axil_arready),   // output wire s_axi_arready
  .probe16(m_axil_rdata),       // output wire [31 : 0] s_axi_rdata
  .probe17(m_axil_rresp),       // output wire [1 : 0] s_axi_rresp
  .probe18(m_axil_rvalid),     // output wire s_axi_rvalid
  .probe19(m_axil_rready),     // input wire s_axi_rready
  .probe20(1'b0), // input wire [0:0]  probe20 
  .probe21(8'b0), // input wire [7:0]  probe21 
  .probe22(1'b0), // input wire [0:0]  probe22 
  .probe23(3'b0), // input wire [2:0]  probe23 
  .probe24(2'b0), // input wire [1:0]  probe24 
  .probe25(4'b0), // input wire [0:0]  probe25 
  .probe26(1'b0), // input wire [0:0]  probe26 
  .probe27(8'b0), // input wire [7:0]  probe27 
  .probe28(3'b0), // input wire [2:0]  probe28 
  .probe29(2'b0), // input wire [1:0]  probe29 
  .probe30(1'b0), // input wire [0:0]  probe30 
  .probe31(4'b0), // input wire [3:0]  probe31 
  .probe32(4'b0), // input wire [3:0]  probe32 
  .probe33(4'b0), // input wire [3:0]  probe33 
  .probe34(4'b0), // input wire [3:0]  probe34 
  .probe35(1'b0), // input wire [0:0]  probe35 
  .probe36(4'b0), // input wire [3:0]  probe36 
  .probe37(4'b0), // input wire [3:0]  probe37 
  .probe38(1'b0), // input wire [0:0]  probe38 
  .probe39(1'b0), // input wire [0:0]  probe39 
  .probe40(1'b0), // input wire [0:0]  probe40 
  .probe41(1'b0), // input wire [0:0]  probe41 
  .probe42(1'b0), // input wire [0:0]  probe42  
  .probe43(1'b0) // input wire [0:0]  probe43
);

endmodule
